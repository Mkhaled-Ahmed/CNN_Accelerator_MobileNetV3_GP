module mem_weights();
    